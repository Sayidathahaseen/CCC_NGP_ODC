-- megafunction wizard: %MAX II oscillator%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altufm_osc 

-- ============================================================
-- File Name: oscillator.vhd
-- Megafunction Name(s):
-- 			altufm_osc
--
-- Simulation Library Files(s):
-- 			maxii
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 9.1 Build 222 10/21/2009 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2009 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--altufm_osc CBX_AUTO_BLACKBOX="ALL" OSC_FREQUENCY=300000 osc oscena
--VERSION_BEGIN 9.1 cbx_altufm_osc 2009:10:21:21:22:16:SJ cbx_maxii 2009:10:21:21:22:16:SJ cbx_mgl 2009:10:21:21:37:49:SJ cbx_stratixii 2009:10:21:21:22:16:SJ cbx_util_mgl 2009:10:21:21:22:16:SJ  VERSION_END

 LIBRARY maxii;
 USE maxii.all;

--synthesis_resources = maxii_ufm 1 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  oscillator_altufm_osc_lv5 IS 
	 PORT 
	 ( 
		 osc	:	OUT  STD_LOGIC;
		 oscena	:	IN  STD_LOGIC
	 ); 
 END oscillator_altufm_osc_lv5;

 ARCHITECTURE RTL OF oscillator_altufm_osc_lv5 IS

	 SIGNAL  wire_gnd	:	STD_LOGIC;
	 SIGNAL  wire_vcc	:	STD_LOGIC;
	 SIGNAL  wire_maxii_ufm_block1_osc	:	STD_LOGIC;
	 COMPONENT  maxii_ufm
	 GENERIC 
	 (
		ADDRESS_WIDTH	:	NATURAL := 9;
		ERASE_TIME	:	NATURAL := 500000000;
		INIT_FILE	:	STRING := "UNUSED";
		OSC_SIM_SETTING	:	NATURAL := 180000;
		PROGRAM_TIME	:	NATURAL := 1600000;
		lpm_type	:	STRING := "maxii_ufm"
	 );
	 PORT
	 ( 
		arclk	:	IN STD_LOGIC := '0';
		ardin	:	IN STD_LOGIC := '0';
		arshft	:	IN STD_LOGIC := '1';
		bgpbusy	:	OUT STD_LOGIC;
		busy	:	OUT STD_LOGIC;
		drclk	:	IN STD_LOGIC := '0';
		drdin	:	IN STD_LOGIC := '0';
		drdout	:	OUT STD_LOGIC;
		drshft	:	IN STD_LOGIC := '1';
		erase	:	IN STD_LOGIC := '0';
		osc	:	OUT STD_LOGIC;
		oscena	:	IN STD_LOGIC := '0';
		program	:	IN STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
 BEGIN

	wire_gnd <= '0';
	wire_vcc <= '1';
	osc <= wire_maxii_ufm_block1_osc;
	maxii_ufm_block1 :  maxii_ufm
	  GENERIC MAP (
		ADDRESS_WIDTH => 9,
		OSC_SIM_SETTING => 300000
	  )
	  PORT MAP ( 
		arclk => wire_gnd,
		ardin => wire_gnd,
		arshft => wire_gnd,
		drclk => wire_gnd,
		drdin => wire_gnd,
		drshft => wire_vcc,
		osc => wire_maxii_ufm_block1_osc,
		oscena => oscena
	  );

 END RTL; --oscillator_altufm_osc_lv5
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY oscillator IS
	PORT
	(
		oscena		: IN STD_LOGIC ;
		osc		: OUT STD_LOGIC 
	);
END oscillator;


ARCHITECTURE RTL OF oscillator IS

	SIGNAL sub_wire0	: STD_LOGIC ;



	COMPONENT oscillator_altufm_osc_lv5
	PORT (
			oscena	: IN STD_LOGIC ;
			osc	: OUT STD_LOGIC 
	);
	END COMPONENT;

BEGIN
	osc    <= sub_wire0;

	oscillator_altufm_osc_lv5_component : oscillator_altufm_osc_lv5
	PORT MAP (
		oscena => oscena,
		osc => sub_wire0
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "MAX II"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_PART STRING ""
-- Retrieval info: PRIVATE: INTERFACE_CHOICE NUMERIC "4"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: VERSION_NUMBER NUMERIC "0"
-- Retrieval info: CONSTANT: OSC_FREQUENCY NUMERIC "300000"
-- Retrieval info: USED_PORT: osc 0 0 0 0 OUTPUT NODEFVAL osc
-- Retrieval info: USED_PORT: oscena 0 0 0 0 INPUT NODEFVAL oscena
-- Retrieval info: CONNECT: @oscena 0 0 0 0 oscena 0 0 0 0
-- Retrieval info: CONNECT: osc 0 0 0 0 @osc 0 0 0 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL oscillator.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL oscillator.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL oscillator.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL oscillator.bsf TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL oscillator_inst.vhd FALSE
-- Retrieval info: LIB_FILE: maxii
